module unary_example(
    a,
    y
);
    input a;
    output y;

    assign y = ~a;

endmodule