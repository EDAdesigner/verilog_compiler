// ���ʽ����ģ��
module expression_test(a, b, c, d, out1, out2, out3);
    input a;
    input b;
    input c;
    input d;
    output out1;
    output out2;
    output out3;
    
    wire temp1;
    wire temp2;
    
    // �򵥸�ֵ
    assign temp1 = a & b;
    
    // ���ӱ��ʽ��ֵ
    assign temp2 = (a & b) | (c & d);
    
    // һԪ�����
    assign out1 = ~temp1;
    
    // �����ŵĸ��ӱ��ʽ
    assign out2 = (a & b) | ~(c ^ d);
    
    // �����������ȼ�����
    assign out3 = a & b | c ^ d & ~(a | b) + c - d;
    
endmodule